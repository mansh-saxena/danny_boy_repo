	// megafunction wizard: %FIFO%
	// GENERATION: STANDARD
	// VERSION: WM1.0
	// MODULE: dcfifo 

	// ============================================================
	// File Name: async_fifo.v
	// Megafunction Name(s):
	// 			dcfifo
	//
	// Simulation Library Files(s):
	// 			altera_mf
	// ============================================================
	// ************************************************************
	// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
	//
	// 20.1.0 Build 711 06/05/2020 SJ Lite Edition
	// ************************************************************


	//Copyright (C) 2020  Intel Corporation. All rights reserved.
	//Your use of Intel Corporation's design tools, logic functions 
	//and other software and tools, and any partner logic 
	//functions, and any output files from any of the foregoing 
	//(including device programming or simulation files), and any 
	//associated documentation or information are expressly subject 
	//to the terms and conditions of the Intel Program License 
	//Subscription Agreement, the Intel Quartus Prime License Agreement,
	//the Intel FPGA IP License Agreement, or other applicable license
	//agreement, including, without limitation, that your use is for
	//the sole purpose of programming logic devices manufactured by
	//Intel and sold by Intel or its authorized distributors.  Please
	//refer to the applicable agreement for further details, at
	//https://fpgasoftware.intel.com/eula.


	// synopsys translate_off
	`timescale 1 ps / 1 ps
	// synopsys translate_on
	module async_fifo (
		aclr,
		data,
		rdclk,
		rdreq,
		wrclk,
		wrreq,
		q,
		rdfull,
		wrfull);

		input	  aclr;
		input	[15:0]  data;
		input	  rdclk;
		input	  rdreq;
		input	  wrclk;
		input	  wrreq;
		output	[15:0]  q;
		output	  rdfull;
		output	  wrfull;
	`ifndef ALTERA_RESERVED_QIS
	// synopsys translate_off
	`endif
		tri0	  aclr;
	`ifndef ALTERA_RESERVED_QIS
	// synopsys translate_on
	`endif

		wire [15:0] sub_wire0;
		wire  sub_wire1;
		wire  sub_wire2;
		wire [15:0] q = sub_wire0[15:0];
		wire  rdfull = sub_wire1;
		wire  wrfull = sub_wire2;

		dcfifo	dcfifo_component (
					.aclr (aclr),
					.data (data),
					.rdclk (rdclk),
					.rdreq (rdreq),
					.wrclk (wrclk),
					.wrreq (wrreq),
					.q (sub_wire0),
					.rdfull (sub_wire1),
					.wrfull (sub_wire2),
					.eccstatus (),
					.rdempty (),
					.rdusedw (),
					.wrempty (),
					.wrusedw ());
		defparam
			dcfifo_component.intended_device_family = "Cyclone IV E",
			dcfifo_component.lpm_hint = "MAXIMUM_DEPTH=1024",
			dcfifo_component.lpm_numwords = 1024,
			dcfifo_component.lpm_showahead = "ON",
			dcfifo_component.lpm_type = "dcfifo",
			dcfifo_component.lpm_width = 16,
			dcfifo_component.lpm_widthu = 10,
			dcfifo_component.overflow_checking = "ON",
			dcfifo_component.rdsync_delaypipe = 4,
			dcfifo_component.read_aclr_synch = "OFF",
			dcfifo_component.underflow_checking = "ON",
			dcfifo_component.use_eab = "ON",
			dcfifo_component.write_aclr_synch = "OFF",
			dcfifo_component.wrsync_delaypipe = 4;

	endmodule
