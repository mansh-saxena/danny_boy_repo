`timescale 1ns/1ns
module low_pass_conv_tb;

    localparam TCLK = 20; // 20ns

    localparam W = 32;
    localparam W_FRAC = 16;

    logic clk = 0;
    dstream #(.N(W)) x ();
    dstream #(.N(W)) y ();

    low_pass_conv #(.W(W), .W_FRAC(W_FRAC)) DUT (.*);

    always #(TCLK/2) clk = ~clk;

    localparam LEN = 100;
    logic [W-1:0] audio_data [0:LEN-1] = '{32'h0064_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0032_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0064_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0032_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000,32'h0000_0000};
    logic [W-1:0] expected [0:LEN-1] = '{32'h00000000,32'h00000000,32'h00000000,32'h000007d0,32'h0000189c,32'h00001f40,32'h00000000,32'hffffa04c,32'hfffef598,32'hfffe0f20,32'hfffd1ee4,32'hfffc74f8,32'hfffc76ec,32'hfffd8e9c,32'h00000c4e,32'h00040934,32'h00095b50,32'h000f95a6,32'h00161778,32'h001c25dc,32'h00210cbe,32'h002442d0,32'h00258096,32'h0024cdae,32'h0022851c,32'h001f33b2,32'h001b6994,32'h0017a840,32'h001449f2,32'h00117e52,32'h000f4dc6,32'h000dadc2,32'h000c8e74,32'h000bf00e,32'h000bec26,32'h000caa94,32'h000e4d22,32'h0010de5c,32'h0014434e,32'h00183382,32'h001c3e78,32'h001fd9e8,32'h00227e46,32'h0023bb12,32'h00235d20,32'h002184dc,32'h001e95e2,32'h001b1a7a,32'h0017a840,32'h0014b946,32'h00129508,32'h0011428e,32'h00108ede,32'h0010197c,32'h000f7922,32'h000e5d8a,32'h000c9e46,32'h000a43ee,32'h0007830c,32'h0004ada8,32'h00021c0a,32'h0000189c,32'hfffecd2a,32'hfffe3b76,32'hfffe3a7c,32'hfffe8f72,32'hffff0790,32'hffff7acc,32'hffffd026,32'h00000000,32'h00000fa0,32'h00000c4e,32'h000003e8,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000,32'h00000000};
    logic start = 0;
    initial begin
        $dumpfile("waveform.vcd");
        $dumpvars();
        y.ready = 1'b0;
        #(TCLK*5);
        y.ready = 1'b1;
        start = 1'b1;
        @(posedge x.valid);
        @(negedge x.valid);
        #(TCLK*5);
        $finish();
    end

    // Input Driver:
    integer i = 0;
    always_ff @(posedge clk) begin
        if (start) begin
            x.data <= audio_data[i];
            i <= i < LEN ? i + 1 : LEN;
            x.valid <= i < LEN ? 1'b1 : 1'b0;
        end
    end

    // Output Check:
    logic [W-1:0] expected_output;
    always_ff @(posedge clk) begin
        if (x.ready != y.ready) $error("x.ready != y.ready");
        expected_output <= expected[i];
        if (start) begin
            $display("expected: %h, actual: %h", expected_output, y.data);
            if (expected_output != y.data) $error("Time %d: Expected value %h but got %h.",$time,expected_output,y.data);
        end
    end
    
endmodule
